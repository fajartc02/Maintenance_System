M 10.1607 64.0254 L 20.1607 64.0254 C 20.1607 64.0254 44.3536 64.0254 61 64.0254 C 76.6107 64.0254 84.675 64.0254
100.8036 64.0254 C 116.9321 64.0254 124.9964 64.0254 141.125 64.0254 C 157.2536 64.0254 165.3179 64.0254 181.4464
64.0254 C 197.575 64.0254 205.6393 64.0254 221.7679 64.0254 C 237.8964 64.0254 245.9607 64.0254 262.0893 64.0254 C
278.2179 64.0254 286.2821 64.0254 302.4107 64.0254 C 318.5393 64.0254 326.6036 64.0254 342.7321 64.0254 C 358.8607
64.0254 366.925 64.0254 383.0536 64.0254 C 399.1821 64.0254 407.2464 64.0254 423.375 64.0254 C 439.5036 64.0254 447.5679
64.0254 463.6964 64.0254 C 479.825 64.0254 487.8893 64.0254 504.0179 64.0254 C 520.1464 64.0254 528.2107 64.0254
544.3393 64.0254 C 560.4679 64.0254 568.5321 64.0254 584.6607 64.0254 C 600.7893 64.0254 608.8536 64.0254 624.9821
64.0254 C 641.1107 64.0254 649.175 64.0254 665.3036 64.0254 C 681.4321 64.0254 689.4964 64.0254 705.625 64.0254 C
721.7536 64.0254 729.8179 64.0254 745.9464 64.0254 C 762.075 64.0254 770.1393 64.0254 786.2679 64.0254 C 802.3964
64.0254 810.4607 64.0254 826.5893 64.0254 C 842.7179 64.0254 850.7821 64.0254 866.9107 64.0254 C 883.0393 64.0254
891.1036 64.0254 907.2321 64.0254 C 923.3607 64.0254 931.425 64.0254 947.5536 64.0254 C 963.6821 64.0254 971.7464
64.0254 987.875 64.0254 C 1004.0036 64.0254 1012.0679 64.0254 1028.1964 64.0254 C 1044.325 64.0254 1052.3893 64.0254
1068.5179 64.0254 C 1084.6464 64.0254 1108.8393 64.0254 1108.8393 64.0254 L 1118.8393 64.0254